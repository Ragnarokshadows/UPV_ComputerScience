* C:\Users\Stephane\Desktop\UPV\TCO\Prac5\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Tue May 29 21:03:19 2018



** Analysis setup **
.tran 1n 120n
.OP 
.LIB "C:\Users\Stephane\Desktop\UPV\TCO\Prac5\Schematic1.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
