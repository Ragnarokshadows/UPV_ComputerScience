* C:\Users\Stephane\Desktop\UPV\TCO\Prac4\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Tue May 29 20:05:20 2018



** Analysis setup **
.DC LIN V_VGS 0V 5V 0.1V 
.OP 
.LIB "C:\Users\Stephane\Desktop\UPV\TCO\Prac4\Schematic1.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
